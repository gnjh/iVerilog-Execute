module simple3_tb;

reg [3:0] A;
reg  D;
wire [3:0] B;
wire [3:0] E;

initial
begin
	$dumpfile("simple3_tb.dump");
	$dumpvars;
	#10 {D,A} = 5'b11111;
	#10 {D,A} = 5'b11110;
	#10 {D,A} = 5'b11101;
	#10 {D,A} = 5'b11100;
	#10 {D,A} = 5'b11011;
	#10 {D,A} = 5'b11010;
	#10 {D,A} = 5'b11001;
	#10 {D,A} = 5'b11000;
	#10 {D,A} = 5'b10111;
	#10 {D,A} = 5'b10110;
	#10 {D,A} = 5'b10101;
	#10 {D,A} = 5'b10100;
	#10 {D,A} = 5'b10011;
	#10 {D,A} = 5'b10010;
	#10 {D,A} = 5'b10001;
	#10 {D,A} = 5'b10000;
	#10 {D,A} = 5'b01111;
	#10 {D,A} = 5'b01110;
	#10 {D,A} = 5'b01101;
	#10 {D,A} = 5'b01100;
	#10 {D,A} = 5'b01011;
	#10 {D,A} = 5'b01010;
	#10 {D,A} = 5'b01001;
	#10 {D,A} = 5'b01000;
	#10 {D,A} = 5'b00111;
	#10 {D,A} = 5'b00110;
	#10 {D,A} = 5'b00101;
	#10 {D,A} = 5'b00100;
	#10 {D,A} = 5'b00011;
	#10 {D,A} = 5'b00010;
	#10 {D,A} = 5'b00001;
	#10 {D,A} = 5'b00000;
	#10 $finish;
end

simple3 s (A,D,B,E);

endmodule